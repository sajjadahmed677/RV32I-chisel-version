* Resistor model "short" defined with a fixed resistance of 0.01 ohms.
.model short r r=0.01
* If "short" is called as a subcircuit, then this needs to be supported, too.
.subckt short 1 2 SUB l=0 w=0
R0 1 2 short
.ends
* For diodes called as a subcircuit
* (backwards compatible with earlier PDK version)
.subckt sky130_fd_pr__diode_pw2nd N P a=0 p=0
D0 N P sky130_fd_pr__diode_pw2nd_05v5 area=a
.ends
* (corresponds to current PDK)
.subckt sky130_fd_pr__diode_pw2nd_05v5 N P area=0
D0 N P sky130_fd_pr__diode_pw2nd_05v5 area=area
.ends
* Resistor model "short" defined with a fixed resistance of 0.01 ohms.
.model short r r=0.01
* If "short" is called as a subcircuit, then this needs to be supported, too.
.subckt short 1 2 SUB l=0 w=0
R0 1 2 short
.ends
* For diodes called as a subcircuit
* (backwards compatible with earlier PDK version)
.subckt sky130_fd_pr__diode_pw2nd N P a=0 p=0
D0 N P sky130_fd_pr__diode_pw2nd_05v5 area=a
.ends
* (corresponds to current PDK)
.subckt sky130_fd_pr__diode_pw2nd_05v5 N P area=0
D0 N P sky130_fd_pr__diode_pw2nd_05v5 area=area
.ends
* Resistor model "short" defined with a fixed resistance of 0.01 ohms.
.model short r r=0.01
* If "short" is called as a subcircuit, then this needs to be supported, too.
.subckt short 1 2 SUB l=0 w=0
R0 1 2 short
.ends
* For diodes called as a subcircuit
* (backwards compatible with earlier PDK version)
.subckt sky130_fd_pr__diode_pw2nd N P a=0 p=0
D0 N P sky130_fd_pr__diode_pw2nd_05v5 area=a
.ends
* (corresponds to current PDK)
.subckt sky130_fd_pr__diode_pw2nd_05v5 N P area=0
D0 N P sky130_fd_pr__diode_pw2nd_05v5 area=area
.ends
* Resistor model "short" defined with a fixed resistance of 0.01 ohms.
.model short r r=0.01
* If "short" is called as a subcircuit, then this needs to be supported, too.
.subckt short 1 2 SUB l=0 w=0
R0 1 2 short
.ends
* For diodes called as a subcircuit
* (backwards compatible with earlier PDK version)
.subckt sky130_fd_pr__diode_pw2nd N P a=0 p=0
D0 N P sky130_fd_pr__diode_pw2nd_05v5 area=a
.ends
* (corresponds to current PDK)
.subckt sky130_fd_pr__diode_pw2nd_05v5 N P area=0
D0 N P sky130_fd_pr__diode_pw2nd_05v5 area=area
.ends
